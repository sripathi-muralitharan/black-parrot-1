
package bp_fe_pkg;

  `include "bsg_defines.v"
  `include "bp_common_fe_be_if.vh"
  `include "bp_fe_defines.vh"
  `include "bp_fe_icache.vh"
  `include "bp_fe_mem_defines.vh"
  `include "bp_fe_icache_tag_info.vh"
  `include "bp_fe_icache_stat_info.vh"

endpackage : bp_fe_pkg
